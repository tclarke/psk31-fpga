//
// Author: tclarke
// Licensed under the GNU Public License (GPL) v3
//


module psk31_top (
        input clk,
        input rst
);

dds_sine #(.

endmodule

